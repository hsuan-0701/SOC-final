/////////////////////////////////
//          8bit CLA           //
/////////////////////////////////

    module CLA_8(
        input  wire        Cin,
        input  wire [7:0]  A,
        input  wire [7:0]  B,
        output wire [8:0]  result
    );
        reg [7:0] G, P, S;
        reg [8:0] C;  

        integer i;
        assign result = {C[8], S};

        always @(*) begin
            C[1] = G[0] | (P[0] & C[0]);
            C[2] = G[1] | (P[1] & G[0]) | (P[1] & P[0] & C[0]);
            C[3] = G[2] | (P[2] & G[1]) | (P[2] & P[1] & G[0]) | (P[2] & P[1] & P[0] & C[0]);
            C[4] = G[3] | (P[3] & G[2]) | (P[3] & P[2] & G[1]) | (P[3] & P[2] & P[1] & G[0]) | (P[3] & P[2] & P[1] & P[0] & C[0]);
            C[5] = G[4] | (P[4] & G[3]) | (P[4] & P[3] & G[2]) | (P[4] & P[3] & P[2] & G[1]) | (P[4] & P[3] & P[2] & P[1] & G[0]) | (P[4] & P[3] & P[2] & P[1] & P[0] & C[0]);
            C[6] = G[5] | (P[5] & G[4]) | (P[5] & P[4] & G[3]) | (P[5] & P[4] & P[3] & G[2]) | (P[5] & P[4] & P[3] & P[2] & G[1]) | (P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & C[0]);
            C[7] = G[6] | (P[6] & G[5]) | (P[6] & P[5] & G[4]) | (P[6] & P[5] & P[4] & G[3]) | (P[6] & P[5] & P[4] & P[3] & G[2]) | (P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & C[0]);
            C[8] = G[7] | (P[7] & G[6]) | (P[7] & P[6] & G[5]) | (P[7] & P[6] & P[5] & G[4]) | (P[7] & P[6] & P[5] & P[4] & G[3]) | (P[7] & P[6] & P[5] & P[4] & P[3] & G[2]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & G[1]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & G[0]) | (P[7] & P[6] & P[5] & P[4] & P[3] & P[2] & P[1] & P[0] & C[0]);
        end

        always @(*)begin
            C[0] = Cin;
        end

        always @(*) begin
            for (i = 0; i < 8; i = i + 1) begin
                G[i] = A[i] & B[i];
                P[i] = A[i] ^ B[i];
            end
        end

        always @(*) begin
            for (i = 0; i < 8; i = i + 1)begin
                S[i] = P[i] ^ C[i];
            end
        end

    endmodule